--------------------------------------------------------------------------------
-- Module Name:    CHROM - behavioral
--
-- Author: Aaron Storey
-- 
-- Description: This module generates the character ROM to store the 
--              pixel data for displaying the various characters
-- 
-- 
-- Dependencies: 
-- 
-- 
-- Assisted by:
--
-- Anthonix the great.
-- 
----------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.numeric_std.all;

entity fontrom is port (
  clk25   : in  std_logic;
  address : in  unsigned(8 downto 0);
  data    : out unsigned(7 downto 0)
  );
end fontrom;

architecture behavioral of fontrom is

  type mem_array is array (0 to 511) of unsigned(7 downto 0);
  constant characters : mem_array := (

    --blank character (0)
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",

    --filled character (1)
    "11111111",
    "11111111",
    "11111111",
    "11111111",
    "11111111",
    "11111111",
    "11111111",
    "11111111",

    -- horizontal line (2)
    "00000000",
    "00000000",
    "00000000",
    "11111111",
    "11111111",
    "00000000",
    "00000000",
    "00000000",

    -- vertical line (3)
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",


    -- top right turn (4)
    "00011000",
    "00011000",
    "00011000",
    "00011111",
    "00011111",
    "00000000",
    "00000000",
    "00000000",

    -- top left turn (5)
    "00011000",
    "00011000",
    "00011000",
    "11111000",
    "11111000",
    "00000000",
    "00000000",
    "00000000",

    -- bottom right turn (6)
    "00000000",
    "00000000",
    "00000000",
    "00011111",
    "00011111",
    "00011000",
    "00011000",
    "00011000",

    -- bottom left turn (7)
    "00000000",
    "00000000",
    "00000000",
    "11111000",
    "11111000",
    "00011000",
    "00011000",
    "00011000",

    -- unused (8)
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",

    -- unused (9)
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",

    -- unused (10)
    "00000000",
    "00000000",
    "00000000",
    "11110000",
    "11110000",
    "00000000",
    "00000000",
    "00000000",

    -- unused (11)
    "00000000",
    "00000000",
    "00000000",
    "00001111",
    "00001111",
    "00000000",
    "00000000",
    "00000000",

    -- top head (12)
    "00011000",
    "00011000",
    "00011000",
    "00111100",
    "00111100",
    "00011000",
    "00000000",
    "00000000",

    -- bottom head (13)
    "00000000",
    "00000000",
    "00011000",
    "00111100",
    "00111100",
    "00011000",
    "00011000",
    "00011000",


    -- left head (14)
    "00000000",
    "00000000",
    "00011000",
    "11111100",
    "11111100",
    "00011000",
    "00000000",
    "00000000",

    -- right head (15)
    "00000000",
    "00000000",
    "00011000",
    "00111111",
    "00111111",
    "00011000",
    "00000000",
    "00000000",

    -- unused (16)
    "00000000",
    "11110000",
    "00010000",
    "00010000",
    "11110000",
    "10000000",
    "10000000",
    "00000000",

    -- unused (17)
    "00000000",
    "11110000",
    "00010000",
    "00010000",
    "11110000",
    "10000000",
    "10000000",
    "00000000",

    -- unused (18)
    "00000000",
    "11110000",
    "00010000",
    "00010000",
    "11110000",
    "10000000",
    "10000000",
    "00000000",

    -- unused (19)
    "00000000",
    "11110000",
    "00010000",
    "00010000",
    "11110000",
    "10000000",
    "10000000",
    "00000000",

    -- unused (20)
    "00000000",
    "11110000",
    "00010000",
    "00010000",
    "11110000",
    "10000000",
    "10000000",
    "00000000",

    -- unused (21)
    "00000000",
    "11110000",
    "00010000",
    "00010000",
    "11110000",
    "10000000",
    "10000000",
    "00000000",

    -- unused (22)
    "00000000",
    "11110000",
    "00010000",
    "00010000",
    "11110000",
    "10000000",
    "10000000",
    "00000000",



    -- unused (23)
    "00000000",
    "11110000",
    "00010000",
    "00010000",
    "11110000",
    "10000000",
    "10000000",
    "00000000",

    -- 0  (24)
    "00111000",
    "01000100",
    "01001100",
    "01010100",
    "01100100",
    "01000100",
    "00111000",
    "00000000",


    -- 1  (25)
    "00010000",
    "00110000",
    "00010000",
    "00010000",
    "00010000",
    "00010000",
    "00111000",
    "00000000",

    -- 2 (26)
    "00111000",
    "01000100",
    "00000100",
    "00001000",
    "00010000",
    "00100000",
    "01111100",
    "00000000",

    -- 3 (27)
    "01111100",
    "00001000",
    "00010000",
    "00001000",
    "00000100",
    "01000100",
    "00111000",
    "00000000",

    -- 4 (28)
    "00001000",
    "00011000",
    "00101000",
    "01001000",
    "01111100",
    "00001000",
    "00001000",
    "00000000",

    -- 5 (29)
    "01111100",
    "01000000",
    "01111000",
    "00000100",
    "00000100",
    "01000100",
    "00111000",
    "00000000",

    -- 6 (30)
    "00011000",
    "00100000",
    "01000000",
    "01111000",
    "01000100",
    "01000100",
    "00111000",
    "00000000",

    -- 7 (31)
    "01111100",
    "00000100",
    "00001000",
    "00010000",
    "00100000",
    "00100000",
    "00100000",
    "00000000",

    -- 8 (32)
    "00111000",
    "01000100",
    "01000100",
    "00111000",
    "01000100",
    "01000100",
    "00111000",
    "00000000",

    -- 9 (33)
    "00111000",
    "01000100",
    "01000100",
    "00111000",
    "00000100",
    "00001000",
    "00110000",
    "00000000",


    -- A (34)
    "00111000",
    "01000100",
    "01000100",
    "01000100",
    "01111100",
    "01000100",
    "01000100",
    "00000000",


    -- B (35)
    "01111000",
    "01000100",
    "01000100",
    "01111000",
    "01000100",
    "01000100",
    "01111000",
    "00000000",


    -- C (36)
    "00111000",
    "01000100",
    "01000000",
    "01000000",
    "01000000",
    "01000100",
    "00111000",
    "00000000",


    -- D (37)
    "01110000",
    "01001000",
    "01000100",
    "01000100",
    "01000100",
    "01001000",
    "01110000",
    "00000000",


    -- E (38)
    "01111100",
    "01000000",
    "01000000",
    "01111000",
    "01000000",
    "01000000",
    "01111100",
    "00000000",


    -- F (39)
    "01111100",
    "01000000",
    "01000000",
    "01111000",
    "01000000",
    "01000000",
    "01000000",
    "00000000",


    -- G (40)
    "00111000",
    "01000100",
    "01000000",
    "01011100",
    "01000100",
    "01000100",
    "00111000",
    "00000000",


    -- H (41)
    "01000100",
    "01000100",
    "01000100",
    "01111100",
    "01000100",
    "01000100",
    "01000100",
    "00000000",


    -- I (42)
    "00111000",
    "00010000",
    "00010000",
    "00010000",
    "00010000",
    "00010000",
    "00111000",
    "00000000",


    -- J (43)
    "00011100",
    "00001000",
    "00001000",
    "00001000",
    "00001000",
    "00101000",
    "00110000",
    "00000000",

    -- K (44)
    "01000100",
    "01001000",
    "01010000",
    "01100000",
    "01010000",
    "01001000",
    "01000100",
    "00000000",

    -- L (45)
    "01000000",
    "01000000",
    "01000000",
    "01000000",
    "01000000",
    "01000000",
    "01111100",
    "00000000",

    -- M (46)
    "01000100",
    "01101100",
    "01010100",
    "01000100",
    "01000100",
    "01000100",
    "01000100",
    "00000000",

    -- N (47)
    "01000100",
    "01000100",
    "01100100",
    "01010100",
    "01001100",
    "01000100",
    "01000100",
    "00000000",

    -- O (48)
    "00111000",
    "01000100",
    "01000100",
    "01000100",
    "01000100",
    "01000100",
    "00111000",
    "00000000",

    -- P (49)
    "01111000",
    "01000100",
    "01000100",
    "01111000",
    "01000000",
    "01000000",
    "01000000",
    "00000000",

    -- Q (50)
    "00111000",
    "01000100",
    "01000100",
    "01000100",
    "01010100",
    "01001000",
    "00110100",
    "00000000",

    -- R (51)
    "01111000",
    "01000100",
    "01000100",
    "01111000",
    "01010000",
    "01001000",
    "01000100",
    "00000000",

    -- S (52)
    "00111100",
    "01000000",
    "01000000",
    "00111000",
    "00000100",
    "00000100",
    "01111000",
    "00000000",

    -- T (53)
    "01111100",
    "00010000",
    "00010000",
    "00010000",
    "00010000",
    "00010000",
    "00010000",
    "00000000",

    -- U (54)
    "01000100",
    "01000100",
    "01000100",
    "01000100",
    "01000100",
    "01000100",
    "00111000",
    "00000000",

    -- V (55)
    "01000100",
    "01000100",
    "01000100",
    "01000100",
    "01000100",
    "00101000",
    "00010000",
    "00000000",

    -- W (56)
    "01000100",
    "01000100",
    "01000100",
    "01010100",
    "01010100",
    "01010100",
    "00101000",
    "00000000",

    -- X (57)
    "01000100",
    "01000100",
    "00101000",
    "00010000",
    "00101000",
    "01000100",
    "01000100",
    "00000000",

    -- Y (58)
    "01000100",
    "01000100",
    "01000100",
    "00101000",
    "00010000",
    "00010000",
    "00010000",
    "00000000",

    -- Z (59)
    "01111100",
    "00000100",
    "00001000",
    "00010000",
    "00100000",
    "01000000",
    "01111100",
    "00000000",



    others => (others => '0')
    );
begin

  process (clk25)
  begin
    if clk25'event and clk25 = '1' then
      data <= characters(to_integer(address));
    end if;
  end process;

end behavioral;

library ieee;
use ieee.STD_LOGIC_1164.all;
use ieee.NUMERIC_STD.all;

package gamelogic_pkg is

  type gamelogic_state_t is (IDLE, CHECK, , HEAD_DATA, HEAD_WRITE, CORNER, TAIL_READ, TAIL_WRITE, SCORE, RESET);

end gamelogic_pkg;

package body gamelogic_pkg is



end gamelogic_pkg;

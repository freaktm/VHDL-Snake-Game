--
-- 
--    This Entity contains an array of data elements representing the fonts and characters 

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.numeric_std.ALL;

entity fontrom is Port ( 
	clk25 : in std_logic;
	address: in unsigned(8 downto 0);
	data: 	out unsigned(7 downto 0)
	);
end fontrom;

architecture behavioral of fontrom is

type mem_array is array (0 to 511) of unsigned(7 downto 0);
constant characters: mem_array := (

  --blank square
	"00000000",
	"00000000",
	"00011000",
	"00111111",
	"00111111",
	"00011000",
	"00000000",
	"00000000",
	
  --border square
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",

	-- horizontal line
	"00000000",
	"00000000",
	"00000000",
	"11111111",
	"11111111",
	"00000000",
	"00000000",
	"00000000",
	
	-- vertical line
	"00011000",
	"00011000",
	"00011000",
	"00011000",
	"00011000",
	"00011000",
	"00011000",
	"00011000",
	
	
	-- top right turn
	"00011000",
	"00011000",
	"00011000",
	"00011111",
	"00011111",
	"00000000",
	"00000000",
	"00000000",
	
	-- top left turn
	"00011000",
	"00011000",
	"00011000",
	"11111000",
	"11111000",
	"00000000",
	"00000000",
	"00000000",
	
	-- bottom right turn
	"00000000",
	"00000000",
	"00000000",
	"00011111",
	"00011111",
	"00011000",
	"00011000",
	"00011000",
	
	-- bottom left turn
	"00000000",
	"00000000",
	"00000000",
	"11111000",
	"11111000",
	"00011000",
	"00011000",
	"00011000",
	
	-- top tail
	"00011000",
	"00011000",
	"00011000",
	"00011000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	
	-- bottom tail
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00011000",
	"00011000",
	"00011000",
	"00011000",
	
	-- left tail
	"00000000",
	"00000000",
	"00000000",
	"11110000",
	"11110000",
	"00000000",
	"00000000",
	"00000000",
	
	-- right tail
	"00000000",
	"00000000",
	"00000000",
	"00001111",
	"00001111",
	"00000000",
	"00000000",
	"00000000",
	
	-- top head
	"00011000",
	"00011000",
	"00011000",
	"00111100",
	"00111100",
	"00011000",
	"00000000",
	"00000000",
	
	-- bottom head
	"00000000",
	"00000000",
	"00011000",
	"00111100",
	"00111100",
	"00011000",
	"00011000",
	"00011000",
	
	
	-- left head
	"00000000",
	"00000000",
	"00011000",
	"11111100",
	"11111100",
	"00011000",
	"00000000",
	"00000000",
	
	-- right head
	"00000000",
	"00000000",
	"00011000",
	"00111111",
	"00111111",
	"00011000",
	"00000000",
	"00000000",
	
	-- smash into vertical line
	"00000000",
	"11110000",
	"00010000",
	"00010000",
	"11110000",
	"10000000",
	"10000000",
	"00000000",
	
	-- smash into horizontal line
	"00000000",
	"11110000",
	"00010000",
	"00010000",
	"11110000",
	"10000000",
	"10000000",
	"00000000",
	
	-- smash into topr corner
	"00000000",
	"11110000",
	"00010000",
	"00010000",
	"11110000",
	"10000000",
	"10000000",
	"00000000",
	
	-- smash into topl corner
	"00000000",
	"11110000",
	"00010000",
	"00010000",
	"11110000",
	"10000000",
	"10000000",
	"00000000",
		
	-- smash into bottomr corner
	"00000000",
	"11110000",
	"00010000",
	"00010000",
	"11110000",
	"10000000",
	"10000000",
	"00000000",
	
	-- smash into bottoml corner
	"00000000",
	"11110000",
	"00010000",
	"00010000",
	"11110000",
	"10000000",
	"10000000",
	"00000000",
	
	-- smash into vert tail
	"00000000",
	"11110000",
	"00010000",
	"00010000",
	"11110000",
	"10000000",
	"10000000",
	"00000000",
	

	
	-- smash into horz tail
	"00000000",
	"11110000",
	"00010000",
	"00010000",
	"11110000",
	"10000000",
	"10000000",
	"00000000",

	-- 0
	"00000000",
	"00111100",
	"01100110",
	"01100110",
	"01100110",
	"01100110",
	"00111100",
	"00000000",
	

	-- 1
	"00000000",
	"00011000",
	"00011000",
	"00011000",
	"00011000",
	"00011000",
	"00011000",
	"00000000",

	-- 2
	"00000000",
	"00111100",
	"00001100",
	"00001100",
	"00111100",
	"00100000",
	"00100000",
	"00000000",

	-- 3
	"00000000",
	"11110000",
	"00010000",
	"00010000",
	"11110000",
	"10000000",
	"10000000",
	"00000000",

	-- 4
	"00000000",
	"11110000",
	"00010000",
	"00010000",
	"11110000",
	"10000000",
	"10000000",
	"00000000",

	-- 5
	"00000000",
	"11110000",
	"00010000",
	"00010000",
	"11110000",
	"10000000",
	"10000000",
	"00000000",

	-- 6
	"00000000",
	"11110000",
	"00010000",
	"00010000",
	"11110000",
	"10000000",
	"10000000",
	"00000000",

	-- 7
	"00000000",
	"11110000",
	"00010000",
	"00010000",
	"11110000",
	"10000000",
	"10000000",
	"00000000",

	-- 8
	"00000000",
	"11110000",
	"00010000",
	"00010000",
	"11110000",
	"10000000",
	"10000000",
	"00000000",

	-- 9
	"00000000",
	"11110000",
	"00010000",
	"00010000",
	"11110000",
	"10000000",
	"10000000",
	"00000000",
	
	
	-- A
	"00000000",
	"11110000",
	"00010000",
	"00010000",
	"11110000",
	"10000000",
	"10000000",
	"00000000",
	
	
	-- B
	"00000000",
	"11110000",
	"00010000",
	"00010000",
	"11110000",
	"10000000",
	"10000000",
	"00000000",
	
	
	-- C
	"00000000",
	"11110000",
	"00010000",
	"00010000",
	"11110000",
	"10000000",
	"10000000",
	"00000000",
	
	
	-- D
	"00000000",
	"11110000",
	"00010000",
	"00010000",
	"11110000",
	"10000000",
	"10000000",
	"00000000",
	
	
	-- E
	"00000000",
	"11110000",
	"00010000",
	"00010000",
	"11110000",
	"10000000",
	"10000000",
	"00000000",
	
	
	-- F
	"00000000",
	"11110000",
	"00010000",
	"00010000",
	"11110000",
	"10000000",
	"10000000",
	"00000000",
	
	
	-- G
	"00000000",
	"11110000",
	"00010000",
	"00010000",
	"11110000",
	"10000000",
	"10000000",
	"00000000",
	
	
	-- H
	"00000000",
	"11110000",
	"00010000",
	"00010000",
	"11110000",
	"10000000",
	"10000000",
	"00000000",
	
	
	-- I
	"00000000",
	"11110000",
	"00010000",
	"00010000",
	"11110000",
	"10000000",
	"10000000",
	"00000000",
	
	
	-- J
	"00000000",
	"11110000",
	"00010000",
	"00010000",
	"11110000",
	"10000000",
	"10000000",
	"00000000",
	
	-- K
	"00000000",
	"11110000",
	"00010000",
	"00010000",
	"11110000",
	"10000000",
	"10000000",
	"00000000",
	
	-- L
	"00000000",
	"11110000",
	"00010000",
	"00010000",
	"11110000",
	"10000000",
	"10000000",
	"00000000",
	
	-- M
	"00000000",
	"11110000",
	"00010000",
	"00010000",
	"11110000",
	"10000000",
	"10000000",
	"00000000",
	
	-- N
	"00000000",
	"11110000",
	"00010000",
	"00010000",
	"11110000",
	"10000000",
	"10000000",
	"00000000",
	
	-- O
	"00000000",
	"11110000",
	"00010000",
	"00010000",
	"11110000",
	"10000000",
	"10000000",
	"00000000",
	
	-- P
	"00000000",
	"11110000",
	"00010000",
	"00010000",
	"11110000",
	"10000000",
	"10000000",
	"00000000",
	
	-- Q
	"00000000",
	"11110000",
	"00010000",
	"00010000",
	"11110000",
	"10000000",
	"10000000",
	"00000000",
	
	-- R
	"00000000",
	"11110000",
	"00010000",
	"00010000",
	"11110000",
	"10000000",
	"10000000",
	"00000000",
	
	-- S
	"00000000",
	"11110000",
	"00010000",
	"00010000",
	"11110000",
	"10000000",
	"10000000",
	"00000000",
	
	-- T
	"00000000",
	"11110000",
	"00010000",
	"00010000",
	"11110000",
	"10000000",
	"10000000",
	"00000000",
	
	-- U
	"00000000",
	"11110000",
	"00010000",
	"00010000",
	"11110000",
	"10000000",
	"10000000",
	"00000000",
	
	-- V
	"00000000",
	"11110000",
	"00010000",
	"00010000",
	"11110000",
	"10000000",
	"10000000",
	"00000000",
	
	-- W
	"00000000",
	"11110000",
	"00010000",
	"00010000",
	"11110000",
	"10000000",
	"10000000",
	"00000000",
	
	-- X
	"00000000",
	"11110000",
	"00010000",
	"00010000",
	"11110000",
	"10000000",
	"10000000",
	"00000000",
	
	-- Y
	"00000000",
	"11110000",
	"00010000",
	"00010000",
	"11110000",
	"10000000",
	"10000000",
	"00000000",
	
	-- Z
	"00000000",
	"11110000",
	"00010000",
	"00010000",
	"11110000",
	"10000000",
	"10000000",
	"00000000",
	

	
	others => (others => '0')
);
begin

process (clk25)
begin
	if clk25'event and clk25='1' then
		data <= characters(to_integer(address));
   end if;
end process;

end behavioral;